* EESchema Netlist Version 1.1 (Spice format) creation date: 4/12/2014 1:56:52 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
K1  N-000005 GND N-000004 15VAC		
BR1  N-000005 N-000004 N-000012 N-000013 2KBP06M-E4/45		
C1  N-000012 N-000003 .47u		
C3  N-000012 GND .47u		
C2  N-000003 N-000013 .47u		
C4  GND N-000013 .47u		
U3  N-000012 GND N-000010 LM7815CT		
U4  GND N-000013 N-000011 LM7915CT		
C8  N-000010 GND 0.1u		
C9  GND N-000011 0.1u		
D3  GND N-000010 1N4001		
D4  N-000011 GND 1N4001		
U2  N-000012 N-000019 GND N-000009 GND LM2596S-ADJ		
R1  N-000012 N-000009 1K		
R2  N-000009 N-000001 6.34K 1%		
D2  GND N-000019 1N5825		
L2  N-000019 N-000001 47u		
C7  N-000001 GND 330u/25V		
C5  N-000009 N-000001 1.5n		
U1  N-000012 N-000014 GND N-000002 GND LM2596SX-3.3		
L1  N-000014 N-000002 37u		
D1  GND N-000014 1N5825		
C6  N-000002 GND 330u/25V		
P1  N-000002 N-000001 N-000010 N-000011 GND GND CONN_6		
C11  ? ? CP1		
C10  ? GND 120u/35V		

.end
